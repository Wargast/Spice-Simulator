entity 
